
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: CQU
// Engineer: Napbad
// 
// Create Date: 12/24/2024 04:23:00 PM
// Design Name: cqu_mips
// Module Name: cache_inst
// Project Name: cqu_mips
// Target Devices: 
// Tool Versions: 
// Description: This cache module implements the instruction cache functionality in the MIPS processor.
//              This module handles read operations of instruction, manages cache coherence, and interacts with the
//              memory and other modules in the datapath.
// 
// Dependencies: 
// - Memory module (mem)
// - Control unit (control)
// - Datapath module (datapath)
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// - This module is part of the MIPS processor design aimed at implementing a complete five-stage pipeline architecture.
// - Ensure that the correct tool versions are used during simulation and synthesis.
// 
//////////////////////////////////////////////////////////////////////////////////
